module top_module (
    input clk,
    input resetn,    // active-low synchronous reset
    input x,
    input y,
    output f,
    output g
); 

    parameter A=4'd0, f1=4'd1, tmp1=4'd2, tmp2=4'd3, g1=4'd4, g1p=4'd5, tmp3=4'd6, g0p=4'd7, tmp0=4'd8;
    reg	[3:0] state, next_state;
    
    always@(*) begin
        case(state)
            A: begin
                if(resetn) 
                    next_state = f1;
                else
                    next_state = A;
            end
            f1:		next_state = tmp0;
            tmp0: begin
                if(x)
                    next_state = tmp1;
                else
                    next_state = g0p;
            end
            tmp1: begin
                if(~x)
                    next_state = tmp2;
                else
                    next_state = g0p;
            end
            tmp2: begin
                if(x)
                    next_state = g1;
                else
                    next_state = g0p;
            end
            g1:	begin
                if(y)
                    next_state = g1p;
                else
                    next_state = tmp3;
            end
            tmp3: begin
                if(y)
                    next_state = g1p;
                else
                    next_state = g0p;
            end
            g1p: begin
                if(~resetn)
                    next_state = A;
                else
                    next_state = g1p;
            end
            g0p: begin
                if(~resetn)
                    next_state = A;
                else
                    next_state = g0p;
            end
        endcase
    end
    
    always@(posedge clk) begin
        if(~resetn)
            state <= A;
        else
            state <= next_state;
    end
    
    assign	f = (state==f1);
    assign	g = (state==g1 || state==tmp3 || state==g1p);
    
endmodule
